<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-32.0494,25.4777,129.982,-65.2201</PageViewport>
<gate>
<ID>2</ID>
<type>AE_RAM_8x8</type>
<position>12.5,-19</position>
<input>
<ID>ADDRESS_0</ID>11 </input>
<input>
<ID>ADDRESS_1</ID>12 </input>
<input>
<ID>ADDRESS_2</ID>7 </input>
<input>
<ID>ADDRESS_3</ID>6 </input>
<input>
<ID>ADDRESS_4</ID>5 </input>
<input>
<ID>ADDRESS_5</ID>4 </input>
<input>
<ID>ADDRESS_6</ID>3 </input>
<input>
<ID>ADDRESS_7</ID>2 </input>
<input>
<ID>DATA_IN_0</ID>19 </input>
<input>
<ID>DATA_IN_1</ID>20 </input>
<input>
<ID>DATA_IN_2</ID>21 </input>
<input>
<ID>DATA_IN_3</ID>22 </input>
<input>
<ID>DATA_IN_4</ID>23 </input>
<input>
<ID>DATA_IN_5</ID>24 </input>
<input>
<ID>DATA_IN_6</ID>26 </input>
<input>
<ID>DATA_IN_7</ID>27 </input>
<output>
<ID>DATA_OUT_0</ID>19 </output>
<output>
<ID>DATA_OUT_1</ID>20 </output>
<output>
<ID>DATA_OUT_2</ID>21 </output>
<output>
<ID>DATA_OUT_3</ID>22 </output>
<output>
<ID>DATA_OUT_4</ID>23 </output>
<output>
<ID>DATA_OUT_5</ID>24 </output>
<output>
<ID>DATA_OUT_6</ID>26 </output>
<output>
<ID>DATA_OUT_7</ID>27 </output>
<input>
<ID>ENABLE_0</ID>18 </input>
<input>
<ID>write_clock</ID>1 </input>
<input>
<ID>write_enable</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 8</lparam>
<lparam>DATA_BITS 8</lparam>
<lparam>Address:0 58</lparam>
<lparam>Address:1 9</lparam>
<lparam>Address:3 198</lparam>
<lparam>Address:4 10</lparam>
<lparam>Address:5 50</lparam>
<lparam>Address:6 10</lparam>
<lparam>Address:8 118</lparam>
<lparam>Address:9 34</lparam>
<lparam>Address:10 44</lparam></gate>
<gate>
<ID>4</ID>
<type>Z-80</type>
<position>34,-23.5</position>
<input>
<ID>/BUSREQ</ID>16 </input>
<output>
<ID>/HALT</ID>31 </output>
<input>
<ID>/INT</ID>31 </input>
<input>
<ID>/NMI</ID>31 </input>
<output>
<ID>/RD</ID>17 </output>
<input>
<ID>/RESET</ID>16 </input>
<input>
<ID>/WAIT</ID>16 </input>
<output>
<ID>/WR</ID>13 </output>
<output>
<ID>A_0</ID>11 </output>
<output>
<ID>A_1</ID>12 </output>
<output>
<ID>A_2</ID>7 </output>
<output>
<ID>A_3</ID>6 </output>
<output>
<ID>A_4</ID>5 </output>
<output>
<ID>A_5</ID>4 </output>
<output>
<ID>A_6</ID>3 </output>
<output>
<ID>A_7</ID>2 </output>
<input>
<ID>CLK</ID>1 </input>
<input>
<ID>D_IN_0</ID>19 </input>
<input>
<ID>D_IN_1</ID>20 </input>
<input>
<ID>D_IN_2</ID>21 </input>
<input>
<ID>D_IN_3</ID>22 </input>
<input>
<ID>D_IN_4</ID>23 </input>
<input>
<ID>D_IN_5</ID>24 </input>
<input>
<ID>D_IN_6</ID>26 </input>
<input>
<ID>D_IN_7</ID>27 </input>
<output>
<ID>D_OUT_0</ID>19 </output>
<output>
<ID>D_OUT_1</ID>20 </output>
<output>
<ID>D_OUT_2</ID>21 </output>
<output>
<ID>D_OUT_3</ID>22 </output>
<output>
<ID>D_OUT_4</ID>23 </output>
<output>
<ID>D_OUT_5</ID>24 </output>
<output>
<ID>D_OUT_6</ID>26 </output>
<output>
<ID>D_OUT_7</ID>27 </output>
<input>
<ID>GND</ID>32 </input>
<input>
<ID>VCC</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>A 2C</lparam>
<lparam>A' </lparam>
<lparam>B </lparam>
<lparam>B' </lparam>
<lparam>C </lparam>
<lparam>C' </lparam>
<lparam>D </lparam>
<lparam>D' </lparam>
<lparam>E </lparam>
<lparam>E' </lparam>
<lparam>F 00</lparam>
<lparam>F' </lparam>
<lparam>H </lparam>
<lparam>H' </lparam>
<lparam>HEX_DISP 000000</lparam>
<lparam>I 00</lparam>
<lparam>IFF1 0</lparam>
<lparam>IFF2 0</lparam>
<lparam>IMF 0</lparam>
<lparam>INFO_STRING opp\3A\20HALT\0A\0Adescription\3A\20Stops\20the\20machine\20until\20it\20is\20reset\20or\20an\20interrupt\20is\20received\0A</lparam>
<lparam>IX </lparam>
<lparam>IY </lparam>
<lparam>L </lparam>
<lparam>L' </lparam>
<lparam>PAUSE_SIM TRUE</lparam>
<lparam>PC 0009</lparam>
<lparam>R 00</lparam>
<lparam>SP </lparam>
<lparam>ZAD_MODE SMART</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_INVERTER</type>
<position>48,-36</position>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8</ID>
<type>EE_VDD</type>
<position>62.5,-30.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_INVERTER</type>
<position>50.5,-40.5</position>
<input>
<ID>IN_0</ID>17 </input>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>12</ID>
<type>EE_VDD</type>
<position>2,-24</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>14</ID>
<type>EE_VDD</type>
<position>-0.5,-34.5</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>18</ID>
<type>FF_GND</type>
<position>49.5,-27.5</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>BB_CLOCK</type>
<position>9.5,9.5</position>
<output>
<ID>CLK</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-17.2,24,-15</points>
<intersection>-17.2 1</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-17.2,25,-17.2</points>
<connection>
<GID>4</GID>
<name>CLK</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-15,24,-15</points>
<intersection>17.5 4</intersection>
<intersection>21 5</intersection>
<intersection>24 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>17.5,-17.5,17.5,-15</points>
<connection>
<GID>2</GID>
<name>write_clock</name></connection>
<intersection>-15 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>21,-15,21,9.5</points>
<intersection>-15 2</intersection>
<intersection>9.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>13.5,9.5,21,9.5</points>
<connection>
<GID>20</GID>
<name>CLK</name></connection>
<intersection>21 5</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-7,25,-6.9</points>
<intersection>-7 1</intersection>
<intersection>-6.9 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7.5,-7,25,-7</points>
<intersection>7.5 3</intersection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-6.9,43,-6.9</points>
<intersection>25 0</intersection>
<intersection>43 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>7.5,-15.5,7.5,-7</points>
<connection>
<GID>2</GID>
<name>ADDRESS_7</name></connection>
<intersection>-7 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>43,-14.4,43,-6.9</points>
<connection>
<GID>4</GID>
<name>A_7</name></connection>
<intersection>-6.9 2</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-15.8,44,-6</points>
<intersection>-15.8 2</intersection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-6,44,-6</points>
<intersection>6.5 3</intersection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43,-15.8,44,-15.8</points>
<connection>
<GID>4</GID>
<name>A_6</name></connection>
<intersection>44 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>6.5,-16.5,6.5,-6</points>
<intersection>-16.5 4</intersection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>6.5,-16.5,7.5,-16.5</points>
<connection>
<GID>2</GID>
<name>ADDRESS_6</name></connection>
<intersection>6.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-17.2,45,-5</points>
<intersection>-17.2 2</intersection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5.5,-5,45,-5</points>
<intersection>5.5 3</intersection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43,-17.2,45,-17.2</points>
<connection>
<GID>4</GID>
<name>A_5</name></connection>
<intersection>45 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>5.5,-17.5,5.5,-5</points>
<intersection>-17.5 4</intersection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>5.5,-17.5,7.5,-17.5</points>
<connection>
<GID>2</GID>
<name>ADDRESS_5</name></connection>
<intersection>5.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-18.6,46,-4</points>
<intersection>-18.6 6</intersection>
<intersection>-4 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>4.5,-4,46,-4</points>
<intersection>4.5 3</intersection>
<intersection>46 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>4.5,-18.5,4.5,-4</points>
<intersection>-18.5 4</intersection>
<intersection>-4 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>4.5,-18.5,7.5,-18.5</points>
<connection>
<GID>2</GID>
<name>ADDRESS_4</name></connection>
<intersection>4.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>43,-18.6,46,-18.6</points>
<connection>
<GID>4</GID>
<name>A_4</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-20,47,-3</points>
<intersection>-20 1</intersection>
<intersection>-3 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-20,47,-20</points>
<connection>
<GID>4</GID>
<name>A_3</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3.5,-3,47,-3</points>
<intersection>3.5 3</intersection>
<intersection>47 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>3.5,-19.5,3.5,-3</points>
<intersection>-19.5 4</intersection>
<intersection>-3 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>3.5,-19.5,7.5,-19.5</points>
<connection>
<GID>2</GID>
<name>ADDRESS_3</name></connection>
<intersection>3.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-20.5,2.5,-1.9</points>
<intersection>-20.5 2</intersection>
<intersection>-1.9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2.5,-1.9,48,-1.9</points>
<intersection>2.5 0</intersection>
<intersection>48 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>2.5,-20.5,7.5,-20.5</points>
<connection>
<GID>2</GID>
<name>ADDRESS_2</name></connection>
<intersection>2.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>48,-21.4,48,-1.9</points>
<intersection>-21.4 4</intersection>
<intersection>-1.9 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>43,-21.4,48,-21.4</points>
<connection>
<GID>4</GID>
<name>A_2</name></connection>
<intersection>48 3</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-24.2,50,0</points>
<intersection>-24.2 1</intersection>
<intersection>0 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-24.2,50,-24.2</points>
<connection>
<GID>4</GID>
<name>A_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>0.5,0,50,0</points>
<intersection>0.5 3</intersection>
<intersection>50 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>0.5,-22.5,0.5,0</points>
<intersection>-22.5 4</intersection>
<intersection>0 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>0.5,-22.5,7.5,-22.5</points>
<connection>
<GID>2</GID>
<name>ADDRESS_0</name></connection>
<intersection>0.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-22.8,49,-1</points>
<intersection>-22.8 1</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-22.8,49,-22.8</points>
<connection>
<GID>4</GID>
<name>A_1</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1.5,-1,49,-1</points>
<intersection>1.5 3</intersection>
<intersection>49 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1.5,-21.5,1.5,-1</points>
<intersection>-21.5 4</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>1.5,-21.5,7.5,-21.5</points>
<connection>
<GID>2</GID>
<name>ADDRESS_1</name></connection>
<intersection>1.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-36,44,-35.4</points>
<intersection>-36 1</intersection>
<intersection>-35.4 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-36,45,-36</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43,-35.4,44,-35.4</points>
<connection>
<GID>4</GID>
<name>/WR</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-36,54,-18.5</points>
<intersection>-36 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-18.5,54,-18.5</points>
<connection>
<GID>2</GID>
<name>write_enable</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-36,54,-36</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-32.5,44,-31.2</points>
<intersection>-32.5 2</intersection>
<intersection>-31.2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-31.2,44,-31.2</points>
<connection>
<GID>4</GID>
<name>/BUSREQ</name></connection>
<intersection>43 4</intersection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>44,-32.5,62.5,-32.5</points>
<intersection>44 0</intersection>
<intersection>62.5 8</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>43,-32.6,43,-29.8</points>
<connection>
<GID>4</GID>
<name>/WAIT</name></connection>
<connection>
<GID>4</GID>
<name>/RESET</name></connection>
<intersection>-31.2 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>62.5,-32.5,62.5,-31.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-32.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-40.5,45,-36.8</points>
<intersection>-40.5 1</intersection>
<intersection>-36.8 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-40.5,47.5,-40.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43,-36.8,45,-36.8</points>
<connection>
<GID>4</GID>
<name>/RD</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-40.5,56.5,-19.5</points>
<intersection>-40.5 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-19.5,56.5,-19.5</points>
<connection>
<GID>2</GID>
<name>ENABLE_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53.5,-40.5,56.5,-40.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-28.4,16,-26</points>
<connection>
<GID>2</GID>
<name>DATA_IN_0</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_0</name></connection>
<intersection>-28.4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,-28.4,25,-28.4</points>
<connection>
<GID>4</GID>
<name>D_OUT_0</name></connection>
<connection>
<GID>4</GID>
<name>D_IN_0</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-29.8,15,-26</points>
<connection>
<GID>2</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>2</GID>
<name>DATA_IN_1</name></connection>
<intersection>-29.8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-29.8,25,-29.8</points>
<connection>
<GID>4</GID>
<name>D_OUT_1</name></connection>
<connection>
<GID>4</GID>
<name>D_IN_1</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-26,14,-25.6</points>
<connection>
<GID>2</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>2</GID>
<name>DATA_IN_2</name></connection>
<intersection>-25.6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14,-25.6,25,-25.6</points>
<connection>
<GID>4</GID>
<name>D_OUT_2</name></connection>
<connection>
<GID>4</GID>
<name>D_IN_2</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-27.5,13,-26</points>
<connection>
<GID>2</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>2</GID>
<name>DATA_IN_3</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-27.5,21.5,-27.5</points>
<intersection>13 0</intersection>
<intersection>21.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>21.5,-27.5,21.5,-20</points>
<intersection>-27.5 1</intersection>
<intersection>-20 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>21.5,-20,25,-20</points>
<connection>
<GID>4</GID>
<name>D_OUT_3</name></connection>
<connection>
<GID>4</GID>
<name>D_IN_3</name></connection>
<intersection>21.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-28.1,12,-26</points>
<connection>
<GID>2</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>2</GID>
<name>DATA_IN_4</name></connection>
<intersection>-28.1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-28.1,22.5,-28.1</points>
<intersection>12 0</intersection>
<intersection>22.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>22.5,-28.1,22.5,-18.6</points>
<intersection>-28.1 1</intersection>
<intersection>-18.6 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>22.5,-18.6,25,-18.6</points>
<connection>
<GID>4</GID>
<name>D_OUT_4</name></connection>
<connection>
<GID>4</GID>
<name>D_IN_4</name></connection>
<intersection>22.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-30.9,11,-26</points>
<connection>
<GID>2</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>2</GID>
<name>DATA_IN_5</name></connection>
<intersection>-30.9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11,-30.9,23,-30.9</points>
<intersection>11 0</intersection>
<intersection>23 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>23,-30.9,23,-21.4</points>
<intersection>-30.9 1</intersection>
<intersection>-21.4 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>23,-21.4,25,-21.4</points>
<connection>
<GID>4</GID>
<name>D_OUT_5</name></connection>
<connection>
<GID>4</GID>
<name>D_IN_5</name></connection>
<intersection>23 3</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-31.5,23.5,-22.8</points>
<intersection>-31.5 1</intersection>
<intersection>-22.8 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-31.5,23.5,-31.5</points>
<intersection>10 4</intersection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>23.5,-22.8,25,-22.8</points>
<connection>
<GID>4</GID>
<name>D_OUT_6</name></connection>
<connection>
<GID>4</GID>
<name>D_IN_6</name></connection>
<intersection>23.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>10,-31.5,10,-26</points>
<connection>
<GID>2</GID>
<name>DATA_IN_6</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_6</name></connection>
<intersection>-31.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-32.5,24,-27</points>
<intersection>-32.5 1</intersection>
<intersection>-27 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-32.5,24,-32.5</points>
<intersection>9 4</intersection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>24,-27,25,-27</points>
<connection>
<GID>4</GID>
<name>D_OUT_7</name></connection>
<connection>
<GID>4</GID>
<name>D_IN_7</name></connection>
<intersection>24 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>9,-32.5,9,-26</points>
<connection>
<GID>2</GID>
<name>DATA_IN_7</name></connection>
<connection>
<GID>2</GID>
<name>DATA_OUT_7</name></connection>
<intersection>-32.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4,-25,4,-24.2</points>
<intersection>-25 2</intersection>
<intersection>-24.2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,-24.2,25,-24.2</points>
<connection>
<GID>4</GID>
<name>VCC</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>2,-25,4,-25</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>4 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-35.5,2,-31.2</points>
<intersection>-35.5 2</intersection>
<intersection>-31.2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-31.2,25,-31.2</points>
<connection>
<GID>4</GID>
<name>/INT</name></connection>
<intersection>2 0</intersection>
<intersection>21.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-0.5,-35.5,2,-35.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>2 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>21.5,-34,21.5,-31.2</points>
<intersection>-34 5</intersection>
<intersection>-32.6 6</intersection>
<intersection>-31.2 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>21.5,-34,25,-34</points>
<connection>
<GID>4</GID>
<name>/HALT</name></connection>
<intersection>21.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>21.5,-32.6,25,-32.6</points>
<connection>
<GID>4</GID>
<name>/NMI</name></connection>
<intersection>21.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-26.5,49.5,-25.6</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>-25.6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-25.6,49.5,-25.6</points>
<connection>
<GID>4</GID>
<name>GND</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,113.8,-63.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,113.8,-63.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,113.8,-63.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,113.8,-63.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,113.8,-63.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,113.8,-63.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,113.8,-63.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,113.8,-63.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,113.8,-63.7</PageViewport></page 9></circuit>